class transaction;
   rand bit[7:0] din;
   rand bit[7:0] addr;
  bit cs;
   bit we;
    bit rd;
  logic clk;
  //bit[7:0] sram_out;
  bit[7:0] dout;
endclass
