module func_return_void;
  
  initial
  begin
    disp("\t passing string to function for displaying");
    disp("\t passing string to function for displaying");
  end

    $display("%s",str);
  endfunction : disp

endmodule : func_return_void
