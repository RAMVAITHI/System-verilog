interface operation;
  logic clk,rst;
  bit [3:0]q;
endinterface
