class transaction;
  logic clk;
  logic rst;
  bit [3:0]q;
endclass
